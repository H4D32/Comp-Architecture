`timescale 1ns/1ps
`include "alu.v"

module alu_test;

    reg[31:0] instruction, reg_A, reg_B;

    wire signed [31:0] result;
    wire[2:0] flags;

    alu test_alu(instruction, reg_A, reg_B,result,flags);

    initial begin

        $display("Format: ");
        $monitor("whole instruction: \n|%32b| \n|opcode|rs(hex) |rt(hex) |\n|%6b|%h|%h| \nfunction(R-types)\n|%6b| \nreg_A(hex)\t: |%h| \nreg_B(hex)\t: |%h| \nresult(hex)\t: |%h| \nflags\t\t: |%3b| \n",
        instruction, test_alu.opcode, test_alu.RSBuffer, test_alu.RTBuffer, test_alu.funct, reg_A, reg_B, result, flags);

        #10 
        $display("Add");
        instruction <= 32'b0000_0000_0010_0000_0101_1000_0010_0000; //add $t3, $reg_B, $reg_A
        reg_A <= 32'b0000_0000_0000_0000_0001_0010_1111_1101; //decimal 4861
        reg_B <= 32'b0000_0000_0000_0000_0001_0110_1111_0010; //decimal 5874

        #10 
        $display("Add (overflow)");
        instruction <= 32'b0000_0000_0010_0000_0101_1000_0010_0000; //add $t3, $reg_B, $reg_A
        reg_A <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
        reg_B <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;        
        
        #10 
        $display("Addu");
        instruction <= 32'b0000_0000_0000_0001_0101_1000_0010_0001; //addu $t3, $reg_A, $reg_B 
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

        #10 
        $display("Sub");
        instruction <= 32'b0000_0000_0000_0001_0000_1000_0010_0010; //sub $at, $reg_A, $reg_B
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0001_0100; //decimal 20
        
        #10 
        $display("Subu");
        instruction <= 32'b0000_0000_0000_0001_1100_1000_0010_0011; //subu $t9, $reg_A, $reg_B
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1001; //decimal 9
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0010; //decimal 2 

        #10
        $display("Addi");
        instruction <= 32'b0010_0000_0000_0000_0000_0010_1011_1100; //addi $zero, $reg_A, 700 
        reg_A <= 32'b0000_0010_0000_0010_0000_0011_1110_1000; // decimal 1000 
        reg_B <= 32'b1000_0000_0000_0010_0000_0000_0001_0001;

        #10 
        $display("Addiu");
        instruction <= 32'b0010_0100_0010_0010_0000_0000_0001_0100; //addiu $v0, $reg_B, 20
        reg_A <= 32'b0000_0000_0000_0000_0000_0001_0000_0000;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

        #10
        $display("And"); 
        instruction <= 32'b0000_0000_0010_0000_0000_0000_0010_0100; //and $zero, $reg_B, $reg_A
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1100; //result should be Reg A
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_1101;

        #10 
        $display("Andi");
        instruction <= 32'b0011_0000_0000_0001_0000_0000_0000_1111; //andi $at, $reg_A, 15
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1100; //result should be Reg A
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

        #10 
        $display("Or");
        instruction <= 32'b0000_0000_0010_0000_1000_0000_0010_0101; //or $s0, $reg_B, $reg_A
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1000; //result 1100 
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;

        #10 
        $display("Nor");
        instruction <= 32'b0000_0000_0000_0001_1001_0000_0010_0111; //nor $s2, $reg_A, $reg_B
        reg_A <= 32'b1111_1111_1111_1111_1111_1111_1111_0001; //result 1100 
        reg_B <= 32'b1111_1111_1111_1111_1111_1111_1111_0010; 

        #10 
        $display("Xor");
        instruction <= 32'b0000_0000_0010_0000_0001_1000_0010_0110; //xor $v1, $reg_B, $reg_A
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1001; //result 1100 
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;

        #10 
        $display("Ori");
        instruction <= 32'b0011_0100_0001_0001_1111_1111_1111_1010; //ori $s1, $reg_A, -6
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0001_0100;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

        #10 
        $display("Xori");
        instruction <= 32'b0011_1000_0010_1111_0000_0000_0000_1100; //xori $t7, $reg_B, 12
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_1001;

        #10 
        $display("Slt");
        instruction <= 32'b0000_0000_0010_0000_0111_0000_0010_1010; //slt $t6, $reg_B, $reg_A
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

        #10 
        $display("Sltu");
        instruction <= 32'b0000_0000_0000_0001_1001_0000_0010_1011; //sltu $s2, $reg_A, $reg_B
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0110;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0001_0001;

        #10 
        $display("Slti");
        instruction <= 32'b0010_1000_0000_1000_1111_1111_1111_1010; //slti $t0, $reg_A, -6
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

        #10 
        $display("Sltiu");
        instruction <= 32'b0010_1100_0010_1011_0000_0000_0000_0100; //sltiu $t3, $reg_B, 4
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        reg_B <= 32'b1111_1111_1111_1111_1111_1111_1111_1010;

        #10 
        $display("Sll");
        instruction <= 32'b0000_0000_0000_0001_0111_1001_0000_0000; //sll $t7, $reg_B, 4
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        reg_B <= 32'b1100_1100_1100_1100_1100_1100_1100_1100; //shift by 4 bits - 1 hexa digit

        #10 
        $display("Sllv");
        instruction <= 32'b0000_0000_0010_0000_1011_1000_0000_0100; //sllv $s7, $reg_A, $reg_B
        reg_A <= 32'b1100_1100_1100_1100_1100_1100_1100_1100;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0100; //shift by 4 bits - 1 hexa digit

        #10 
        $display("Srl");
        instruction <= 32'b0000_0000_0000_0000_0111_0001_0000_0010; //srl $t6, $reg_A, 4
        reg_A <= 32'b1100_1100_1100_1100_1100_1100_1100_1100;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0100; //shift by 4 bits - 1 hexa digit

        #10 
        $display("Srlv");
        instruction <= 32'b0000_0000_0000_0001_1100_1000_0000_0110; //srlv $t9, $reg_B, $reg_A
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0100; //shift by 4 bits - 1 hexa digit
        reg_B <= 32'b1100_1100_1100_1100_1100_1100_1100_1100;

        #10 
        $display("Sra");
        instruction <= 32'b0000_0000_0000_0000_0101_1001_0000_0011; //sra $t3, $reg_A, 4
        reg_A <= 32'b1100_1100_1100_1100_1100_1100_1100_1100;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

        #10 
        $display("Srav");
        instruction <= 32'b0000_0000_0010_0000_0000_0000_0000_0111; //srav $s8, $reg_A, $reg_B
        reg_A <= 32'b1100_1100_1100_1100_1100_1100_1100_1100;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;

        #10 
        $display("Beq - Success");
        instruction <= 32'b0001_0000_0010_0000_0000_0000_0000_1100; //beq $reg_B, $reg_A, 12
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

        #10 
        $display("Bne - Fail");
        instruction <= 32'b0001_0100_0000_0001_0000_0000_0000_1100; //bne $reg_A, $reg_B, 12
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

        #10 
        $display("Lw");
        instruction <= 32'b1000_1100_0011_0000_0000_0000_0000_0000; //lw $s0, 0($reg_B)
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        reg_B <= 32'b0000_0000_0000_0000_0000_1000_0001_0000;

        #10 
        $display("Sw");
        instruction <= 32'b1010_1100_0000_1000_0000_0000_0000_1000; //sw $t0, 8($reg_A)
        reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
        
        #10 $finish;
    end
endmodule